module top(
);

endmodule : top
