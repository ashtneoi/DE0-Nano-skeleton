module test(
);

endmodule : test
